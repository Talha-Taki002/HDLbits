module top_module(output wire out, input wire in);
    assign out = ~in;
endmodule