module top_module(input wire a, b, c, output wire w, x, y, z);
    assign w = a, x = b, y = b, z = c;
endmodule