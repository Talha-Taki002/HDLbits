module top_module(output out, input a, b);
    assign out = ~ (a | b);
endmodule