module top_module(output wire out, input wire a, b);
    assign out = a & b;
endmodule